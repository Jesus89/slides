module led(output wire LED);
  assign LED = 1'b1;
endmodule
